/////////////////////////////////////////////////////////////////////////////////////
// File Name : axi.svh
// Version   : 0.1
//-------------------axi.svh------------------------------------
/////////////////////////////////////////////////////////////////////////////////////

    
`ifndef AXI_SVH
`define AXI_SVH

  `include "axi_packet.sv"
  `include "axi_monitor.sv"
  `include "axi_sequencer.sv"	
  `include "axi_sequence.sv"
  `include "axi_driver.sv"
  `include "axi_agent.sv"
  `include "axi_scoreboard.sv"
  `include "axi_env.sv"
 
`endif// AXI_SVH


